// Copyright (C) 2020  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// Generated by Quartus Prime Version 20.1.1 Build 720 11/11/2020 SJ Lite Edition
// Created on Wed Dec 22 20:41:43 2021

// synthesis message_off 10175

`timescale 1ns/1ns

module control_unit (
    reset,clock,dipor,cnt,dip8,
    player,progress,terminate);

    input reset;
    input clock;
    input dipor;
    input [1:0] cnt;
    input dip8;
    tri0 reset;
    tri0 dipor;
    tri0 [1:0] cnt;
    tri0 dip8;
    output player;
    output progress;
    output terminate;
    reg player;
    reg progress;
    reg terminate;
    reg [6:0] fstate;
    reg [6:0] reg_fstate;
    parameter state1=0,state3=1,state2=2,state5=3,state6=4,state4=5,state7=6;

    always @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
        end
    end

    always @(fstate or reset or dipor or cnt or dip8)
    begin
        if (~reset) begin
            reg_fstate <= state1;
            player <= 1'b0;
            progress <= 1'b0;
            terminate <= 1'b0;
        end
        else begin
            player <= 1'b0;
            progress <= 1'b0;
            terminate <= 1'b0;
            case (fstate)
                state1: begin
                    if (((dipor == 1'b1) & (dip8 == 1'b1)))
                        reg_fstate <= state1;
                    else if (((dipor == 1'b0) & (dip8 == 1'b1)))
                        reg_fstate <= state2;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state1;

                    player <= 1'b0;

                    progress <= 1'b0;

                    terminate <= 1'b0;
                end
                state3: begin
                    if (((dipor == 1'b1) & (dip8 == 1'b1)))
                        reg_fstate <= state4;
                    else if ((dip8 == 1'b0))
                        reg_fstate <= state1;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state3;

                    player <= 1'b1;

                    progress <= 1'b1;

                    terminate <= 1'b0;
                end
                state2: begin
                    if (((dipor == 1'b0) & (dip8 == 1'b1)))
                        reg_fstate <= state2;
                    else if (((dipor == 1'b1) & (dip8 == 1'b1)))
                        reg_fstate <= state3;
                    else if ((dip8 == 1'b0))
                        reg_fstate <= state1;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state2;

                    player <= 1'b1;

                    progress <= 1'b0;

                    terminate <= 1'b0;
                end
                state5: begin
                    if (((dipor == 1'b0) & (dip8 == 1'b1)))
                        reg_fstate <= state5;
                    else if (((dipor == 1'b1) & (dip8 == 1'b1)))
                        reg_fstate <= state6;
                    else if ((dip8 == 1'b0))
                        reg_fstate <= state1;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state5;

                    player <= 1'b0;

                    progress <= 1'b0;

                    terminate <= 1'b0;
                end
                state6: begin
                    if (((cnt[1:0] != 2'b10) | (dip8 == 1'b0)))
                        reg_fstate <= state1;
                    else if (((cnt[1:0] == 2'b10) & (dip8 == 1'b1)))
                        reg_fstate <= state7;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state6;

                    player <= 1'b0;

                    progress <= 1'b1;

                    terminate <= 1'b0;
                end
                state4: begin
                    if (((dipor == 1'b0) & (dip8 == 1'b1)))
                        reg_fstate <= state5;
                    else if (((dipor == 1'b1) & (dip8 == 1'b1)))
                        reg_fstate <= state4;
                    else if ((dip8 == 1'b0))
                        reg_fstate <= state1;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state4;

                    player <= 1'b1;

                    progress <= 1'b0;

                    terminate <= 1'b0;
                end
                state7: begin
                    if (((cnt[1:0] == 2'b10) & (dip8 == 1'b1)))
                        reg_fstate <= state7;
                    else if ((dip8 == 1'b0))
                        reg_fstate <= state1;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state7;

                    player <= 1'b0;

                    progress <= 1'b0;

                    terminate <= 1'b1;
                end
                default: begin
                    player <= 1'bx;
                    progress <= 1'bx;
                    terminate <= 1'bx;
                    $display ("Reach undefined state");
                end
            endcase
        end
    end
endmodule // control_unit
