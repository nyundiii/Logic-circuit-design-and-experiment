// Copyright (C) 2020  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// Generated by Quartus Prime Version 20.1.1 Build 720 11/11/2020 SJ Lite Edition
// Created on Wed Dec 08 18:27:42 2021

// synthesis message_off 10175

`timescale 1ns/1ns

module con4 (
    reset,clock,random,trigger,final3,final1,final2,
    final4,En);

    input reset;
    input clock;
    input [3:0] random;
    input trigger;
    input [3:0] final3;
    input [3:0] final1;
    input [3:0] final2;
    tri reset;
    tri [3:0] random;
    tri trigger;
    tri [3:0] final3;
    tri [3:0] final1;
    tri [3:0] final2;
    output [3:0] final4;
    output En;
	 reg [3:0] temprandom;
    reg [3:0] final4;
    reg En;
    reg [4:0] fstate;
    reg [4:0] reg_fstate;
    parameter state1=0,state2=1,state3=2,state4=3;

    always @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
        end
    end

    always @(fstate or reset or random or trigger or final3 or final1 or final2)
    begin
        if (~reset) begin
            reg_fstate <= state1;
            final4 <= 4'b0000;
            En <= 1'b0;
        end
        else begin
            final4 <= 4'b0000;
            En <= 1'b0;
            case (fstate)
                state1: begin
                    if (((trigger == 1'b0) | (final3[3:0] == 4'b0000)))
                        reg_fstate <= state1;
                    else if (((trigger == 1'b1) & (final3[3:0] != 4'b0000)))
                        reg_fstate <= state2;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state1;

                    final4 <= 4'b0000;

                    En <= 1'b0;
                end
                state2: begin
                    if (((((random[3:0] >= 4'b1011) | (random[3:0] == final1[3:0])) | (random[3:0] == final2[3:0])) | (random[3:0] == final3[3:0]))) begin
								
                        reg_fstate <= state2;
								end
                    else if (((((random[3:0] < 4'b1011) & (random[3:0] != final1[3:0])) & (random[3:0] != final2[3:0])) & (random[3:0] != final3[3:0])))
                        reg_fstate <= state3;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state2;

                    final4 <= random[3:0];

                    En <= 1'b1;
                end
                state3: begin
                    if ((final3[3:0] != 4'b0000))
                        reg_fstate <= state4;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state3;

                    final4 <= 4'b0000;

                    En <= 1'b0;
                end
                state4: begin
                    if ((final3[3:0] != 4'b0000))
                        reg_fstate <= state4;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state4;

                    final4 <= 4'b0000;

                    En <= 1'b0;
                end
                
                default: begin
                    final4 <= 4'bxxxx;
                    En <= 1'bx;
                    $display ("Reach undefined state");
                end
            endcase
        end
    end
endmodule // con4
