// Copyright (C) 2020  Intel Corporation. All rights reserved.

// Your use of Intel Corporation's design tools, logic functions 

// and other software and tools, and any partner logic 

// functions, and any output files from any of the foregoing 

// (including device programming or simulation files), and any 

// associated documentation or information are expressly subject 

// to the terms and conditions of the Intel Program License 

// Subscription Agreement, the Intel Quartus Prime License Agreement,

// the Intel FPGA IP License Agreement, or other applicable license

// agreement, including, without limitation, that your use is for

// the sole purpose of programming logic devices manufactured by

// Intel and sold by Intel or its authorized distributors.  Please

// refer to the applicable agreement for further details, at

// https://fpgasoftware.intel.com/eula.

 

// Generated by Quartus Prime Version 20.1.1 Build 720 11/11/2020 SJ Lite Edition

// Created on Thu Dec 09 11:04:54 2021

 

// synthesis message_off 10175

 

`timescale 1ns/1ns

 

module adderpractice (

    reset,clock,inputsum,

    outputsum,carry,ce);

 

    input reset;

    input clock;

    input [4:0] inputsum;

    tri0 reset;

    tri0 [4:0] inputsum;

    output [4:0] outputsum;

	 output carry;

    output ce;

	 reg [4:0] outputsum;

	 reg ce;

	 reg carry;

    reg [4:0] fstate;

    reg [4:0] reg_fstate;

    parameter state1=0,state2=1,state3=2,state4=3,state5=4,state6=5,state7=6,state8=7,state9=8,state10=9,state11=10;

 

    always @(posedge clock)

    begin

        if (clock) begin

            fstate <= reg_fstate;

        end

    end

 

    always @(fstate or reset or inputsum)

    begin

        if (~reset) begin

            reg_fstate <= state1;

            outputsum <= 5'b0_0000;

				carry <= 1'b0;

				ce <= 1'b0;

        end

        else begin

            outputsum <= 5'b0_0000;

				carry <= 1'b0;

				ce <= 1'b0;

            case (fstate)

                state1: begin

                    if ((inputsum[4:0] == 5'b0_1010))

                        reg_fstate <= state2;

                    else if ((inputsum[4:0] == 5'b01011))

                        reg_fstate <= state3;

							else if ((inputsum[4:0] == 5'b01100))

                        reg_fstate <= state4;

							else if ((inputsum[4:0] == 5'b01101))

                        reg_fstate <= state5;

							else if ((inputsum[4:0] == 5'b01110))

                        reg_fstate <= state6;

							else if ((inputsum[4:0] == 5'b01111))

                        reg_fstate <= state7;

							else if ((inputsum[4:0] == 5'b10000))

                        reg_fstate <= state8;

							else if ((inputsum[4:0] == 5'b10001))

                        reg_fstate <= state9;

							else if ((inputsum[4:0] == 5'b10010))

                        reg_fstate <= state10;

							else if ((inputsum[4:0] == 5'b00000))

                        reg_fstate <= state11;
							else
							
								reg_fstate <= state1;

                    // Inserting 'else' block to prevent latch inference

 

                    outputsum <= inputsum[4:0];

						  carry <= 1'b0;

						  ce <= 1'b1;

                end

                state2: begin

		

							reg_fstate <= state1;

 

                    outputsum <= 5'b00000;

						  carry <= 1'b1;

						  ce <= 1'b1;

                end

                state3: begin

                   

                    reg_fstate <= state1;

 

                    outputsum <= 5'b00001;

						  carry <= 1'b1;

						  ce <= 1'b1;

                end

                state4: begin

                    

                    reg_fstate <= state1;

						  ce <= 1'b1;

 

                    outputsum <= 5'b00010;

						  carry <= 1'b1;

                end

					 state5: begin

                    

                    reg_fstate <= state1;

						  ce <= 1'b1;

 

                    outputsum <= 5'b00011;

						  carry <= 1'b1;

                end

					 state6: begin

                    

                    reg_fstate <= state1;

						  ce <= 1'b1;

 

                    outputsum <= 5'b00100;

						  carry <= 1'b1;

                end

					 state7: begin

                    

                    reg_fstate <= state1;

						  ce <= 1'b1;

 

                    outputsum <= 5'b00101;

						  carry <= 1'b1;

                end

					 state8: begin

                    

                    reg_fstate <= state1;

						  ce <= 1'b1;

 

                    outputsum <= 5'b00110;

						  carry <= 1'b1;

                end

					 state9: begin

                    

                    reg_fstate <= state1;

						  ce <= 1'b1;

 

                    outputsum <= 5'b00111;

						  carry <= 1'b1;

                end

					 state10: begin

                    

                    reg_fstate <= state1;

						  ce <= 1'b1;

 

                    outputsum <= 5'b01000;

						  carry <= 1'b1;

                end

					 state11: begin

                    

                    reg_fstate <= state1;

						  ce <= 1'b0;

 

                    outputsum <= 5'b00000;

						  carry <= 1'b0;

                end

                default: begin

                    outputsum <= 5'b00000;

						  carry <= 1'b0;

						  ce <= 1'b0;

                    $display ("Reach undefined state");

                end

            endcase

        end

    end

endmodule // adderpractice