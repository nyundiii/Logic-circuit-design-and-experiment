// Copyright (C) 2020  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// Generated by Quartus Prime Version 20.1.1 Build 720 11/11/2020 SJ Lite Edition
// Created on Wed Dec 22 01:43:26 2021

// synthesis message_off 10175

`timescale 1ns/1ns

module rnd2_ledcontrol (
    reset,clock,inputten,
    ledstate);

    input reset;
    input clock;
    input [3:0] inputten;
    tri reset;
    tri [3:0] inputten;
    output [3:0] ledstate;
    reg [3:0] ledstate;
    reg [4:0] fstate;
    reg [4:0] reg_fstate;
    parameter state1=0,state2=1,state3=2,state4=3,state5=4;

    always @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
        end
    end

    always @(fstate or reset or inputten)
    begin
        if (~reset) begin
            reg_fstate <= state1;
            ledstate <= 4'b0000;
        end
        else begin
            ledstate <= 4'b0000;
            case (fstate)
                state1: begin
                    if (((inputten[3:0] >= 4'b0010) & (inputten[3:0] < 4'b0100)))
                        reg_fstate <= state2;
                    else if (((inputten[3:0] >= 4'b0100) & (inputten[3:0] < 4'b0110)))
                        reg_fstate <= state3;
                    else if (((inputten[3:0] >= 4'b0110) & (inputten[3:0] < 4'b1000)))
                        reg_fstate <= state4;
                    else if ((inputten[3:0] >= 4'b1000))
                        reg_fstate <= state5;
                    else if ((inputten[3:0] < 4'b0010))
                        reg_fstate <= state1;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state1;

                    ledstate <= 4'b1111;
                end
                state2: begin
                    if (((inputten[3:0] >= 4'b0010) & (inputten[3:0] < 4'b0100)))
                        reg_fstate <= state2;
                    else if (((inputten[3:0] >= 4'b0100) & (inputten[3:0] < 4'b0110)))
                        reg_fstate <= state3;
                    else if (((inputten[3:0] >= 4'b0110) & (inputten[3:0] < 4'b1000)))
                        reg_fstate <= state4;
                    else if ((inputten[3:0] >= 4'b1000))
                        reg_fstate <= state5;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state2;

                    ledstate <= 4'b1110;
                end
                state3: begin
                    if (((inputten[3:0] >= 4'b0100) & (inputten[3:0] < 4'b0110)))
                        reg_fstate <= state3;
                    else if (((inputten[3:0] >= 4'b0110) & (inputten[3:0] < 4'b1000)))
                        reg_fstate <= state4;
                    else if ((inputten[3:0] >= 4'b1000))
                        reg_fstate <= state5;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state3;

                    ledstate <= 4'b1100;
                end
                state4: begin
                    if (((inputten[3:0] >= 4'b0110) & (inputten[3:0] < 4'b1000)))
                        reg_fstate <= state4;
                    else if ((inputten[3:0] >= 4'b1000))
                        reg_fstate <= state5;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state4;

                    ledstate <= 4'b1000;
                end
                state5: begin
                    if ((inputten[3:0] >= 4'b1000))
                        reg_fstate <= state5;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state5;

                    ledstate <= 4'b0000;
                end
                default: begin
                    ledstate <= 4'bxxxx;
                    $display ("Reach undefined state");
                end
            endcase
        end
    end
endmodule // rnd2_ledcontrol
