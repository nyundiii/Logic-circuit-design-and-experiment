// Copyright (C) 2020  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// Generated by Quartus Prime Version 20.1.1 Build 720 11/11/2020 SJ Lite Edition
// Created on Tue Dec 21 15:49:51 2021

// synthesis message_off 10175

`timescale 1ns/1ns

module add_b_or_zero (
    reset,clock,reg_out[3:0],ce,
    add_B[3:0]);

    input reset;
    input clock;
    input [3:0] reg_out;
    input ce;
    tri0 reset;
    tri0 [3:0] reg_out;
    tri0 ce;
    output [3:0] add_B;
    reg [3:0] add_B;
    reg [1:0] fstate;
    reg [1:0] reg_fstate;
    parameter state1=0,state2=1;

    always @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
        end
    end

    always @(fstate or reset or reg_out or ce)
    begin
        if (~reset) begin
            reg_fstate <= state1;
            add_B <= 4'b0000;
        end
        else begin
            add_B <= 4'b0000;
            case (fstate)
                state1: begin
                    if ((ce == 1'b0))
                        reg_fstate <= state1;
                    else if ((ce == 1'b1))
                        reg_fstate <= state2;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state1;

                    add_B <= 4'b0000;
                end
                state2: begin
                    reg_fstate <= state1;

                    add_B <= reg_out[3:0];
                end
                default: begin
                    add_B <= 4'bxxxx;
                    $display ("Reach undefined state");
                end
            endcase
        end
    end
endmodule // add_b_or_zero
