// Copyright (C) 2020  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// Generated by Quartus Prime Version 20.1.1 Build 720 11/11/2020 SJ Lite Edition
// Created on Wed Dec 08 23:14:48 2021

// synthesis message_off 10175

`timescale 1ns/1ns

module SBO (
    reset,clock,random,key1,key2,key3,key4,sharp,
    S,B,ce);

    input reset;
    input clock;
    input [3:0] random;
    input [3:0] key1;
	 input [3:0] key2;
	 input [3:0] key3;
	 input [3:0] key4;
    input sharp;
    tri reset;
    tri [3:0] random;
    tri [3:0] key1;
	 tri [3:0] key2;
	 tri [3:0] key3;
	 tri [3:0] key4;
    tri sharp;
    output S;
    output B;
    output ce;
    reg S;
    reg B;
    reg ce;
    reg [4:0] fstate;
    reg [4:0] reg_fstate;
    parameter state2=0,state1=1,state3=2,state4=3,state5=4;

    always @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
        end
    end

    always @(fstate or reset or random or key1 or sharp)
    begin
        if (~reset) begin
            reg_fstate <= state1;
            S <= 1'b0;
            B <= 1'b0;
            ce <= 1'b0;
        end
        else begin
            S <= 1'b0;
            B <= 1'b0;
            ce <= 1'b0;
            case (fstate)
                state2: begin
                    if ((random[3:0] == key1[3:0]))
                        reg_fstate <= state3;
                    else if ((((random[3:0] == key2[3:0]) | (random[3:0] == key3[3:0])) | (random[3:0] == key4[3:0])))
                        reg_fstate <= state4;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state5;

                    S <= 1'b0;

                    B <= 1'b0;

                    ce <= 1'b0;
                end
                state1: begin
                    if ((sharp == 1'b1))
                        reg_fstate <= state2;
                    else if ((sharp == 1'b0))
                        reg_fstate <= state1;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state1;

                    S <= 1'b0;

                    B <= 1'b0;

                    ce <= 1'b0;
                end
                state3: begin
                  
                    reg_fstate <= state1;
                    

                    S <= 1'b1;

                    B <= 1'b0;

                    ce <= 1'b1;
                end
                state4: begin
                    reg_fstate <= state1;
                    

                    S <= 1'b0;

                    B <= 1'b1;

                    ce <= 1'b1;
                end
                state5: begin
                    reg_fstate <= state1;

                    S <= 1'b0;

                    B <= 1'b0;

                    ce <= 1'b1;
                end
                default: begin
                    S <= 1'bx;
                    B <= 1'bx;
                    ce <= 1'bx;
                    $display ("Reach undefined state");
                end
            endcase
        end
    end
endmodule // SBO
